// Emmett Stralka estralka@hmc.edu
// 09/03/25
// Testbench for Lab2_ES module



module Lab2_ES_tb();
    logic clk, reset;
    logic [3:0] s0, s1;
    logic [6:0] seg, seg_expected;
    logic [4:0] led, led_expected;
    logic select;
    logic [31:0] vectornum, errors;
    logic [32:0] testvectors[10000:0]; // Size for: s0(4) + s1(4) + seg_expected(7) + select(1) + led(5) + led_expected(5) = 26 bits

    // Instantiate device under test
    Lab2_ES dut(
        clk,
        s0,
        s1,
        seg,
        led,
        select
    );
    
    // Generate clock (12 MHz - same as main design input clock)
    always begin
        clk = 1; #41.67; clk = 0; #41.67; // 12 MHz = 83.33ns period, 41.67ns half period
    end

    // Clock divider to match the 100 Hz select signal rate
    localparam int HALF_PERIOD = 60_000; // Same as main design
    logic [23:0] divcnt = 0;
    logic test_clk = 0;

    always_ff @(posedge clk) begin
        if (divcnt == HALF_PERIOD - 1) begin
            divcnt <= 0;
            test_clk <= ~test_clk; // 100 Hz test clock
        end else begin
            divcnt <= divcnt + 1;
        end
    end
    
    // Load test vectors and initialize
    initial begin
        $readmemb("Lab2_ES_tb.tv", testvectors);
        vectornum = 0; errors = 0;
        reset = 1; #22; reset = 0;
    end
    
    // Apply test vectors on rising edge of 100 Hz test clock
    always @(posedge test_clk) begin
        if (!reset) begin
            // Test vector format: {s0[3:0], s1[3:0], seg_expected[6:0], select, led[4:0], led_expected[4:0]}
            {s0, s1, seg_expected, select, led, led_expected} = testvectors[vectornum];
        end
    end
    
    // Check results on falling edge of 100 Hz test clock
    always @(negedge test_clk) begin
        if (~reset) begin
            // Check LED output
            if (led !== led_expected) begin
                $display("Error at vector %0d: s0=%b s1=%b | led out %b expected %b", 
                          vectornum, s0, s1, led, led_expected);
                errors = errors + 1;
            end
            
            // Check seven-segment output (multiplexed)
            if (seg !== seg_expected) begin
                $display("Error at vector %0d: s0=%b s1=%b select=%b | seg out %b expected %b", 
                          vectornum, s0, s1, select, seg, seg_expected);
                errors = errors + 1;
            end
            
            vectornum = vectornum + 1;
            if (testvectors[vectornum] === 33'bx) begin
                $display("%d tests completed with %d errors", vectornum, errors);
                $stop;
            end
        end
    end
endmodule
