// Emmett Stralka estralka@hmc.edu
// 09/03/25
// Lab2_ES: Main module implementing a dual seven-segment display system with power multiplexing
module Lab2_ES (
    input  logic        reset,    // Active-low reset signal
    input  logic [3:0]  s0,       // First 4-bit input number
    input  logic [3:0]  s1,       // Second 4-bit input number
    output logic [6:0]  seg,      // Multiplexed seven-segment signal
    output logic [4:0]  led,      // LEDs show sum of s0 + s1
    output logic        select0,  // Power multiplexing control for display 0 (PNP transistor)
    output logic        select1   // Power multiplexing control for display 1 (PNP transistor)
);

    // Clock signal generated by internal oscillator
    logic clk;
    // Internal high-speed oscillator (12 MHz with division factor of 2)
    HSOSC #(.CLKHF_DIV(2'b01)) 
          hf_osc (
              .CLKHFPU(1'b1),  // Power up the oscillator
              .CLKHFEN(1'b1),  // Enable the oscillator
              .CLKHF(clk)      // Output clock signal
          );

    // Internal signals
    logic [4:0] sum;                    // 5-bit sum from adder (s0 + s1)
    logic [6:0] seg0_internal, seg1_internal;  // Seven-segment patterns for each display
    logic display_select;               // Current display selection (0 or 1)
    logic [23:0] divcnt;                // Clock divider counter for multiplexing

    // Seven-segment display decoders for each input number
    seven_segment seven_segment0 (
        .num(s0),              // Input: first 4-bit number
        .seg(seg0_internal)    // Output: 7-segment pattern for s0
    );
    seven_segment seven_segment1 (
        .num(s1),              // Input: second 4-bit number
        .seg(seg1_internal)    // Output: 7-segment pattern for s1
    );

    // 2-to-1 multiplexer for time-multiplexing the seven-segment displays
    MUX2 signal_mux (
        .d0(seg0_internal),    // Input: seven-segment pattern for s0
        .d1(seg1_internal),    // Input: seven-segment pattern for s1
        .select(display_select), // Select signal (0 = s0, 1 = s1)
        .y(seg)                // Output: multiplexed seven-segment signal
    );

    // Five-bit adder to compute sum for LED display
    five_bit_adder adder(
        .s1(s0),    // First 4-bit input
        .s2(s1),    // Second 4-bit input
        .sum(sum)   // 5-bit sum output (handles carry)
    );

    // Output assignments
    assign led = sum;      // LEDs display the sum of s0 + s1 (5 bits)

    // --- Power Multiplexing at ~100 Hz ---
    // This controls which display is powered on to create the illusion of both being on
    localparam int HALF_PERIOD = 60_000; // Half period for 12 MHz input clock (100 Hz switching)

    // Clock divider for power multiplexing
    always_ff @(posedge clk or negedge reset) begin
        if (~reset) begin                    // Async active-low reset
            divcnt <= 0;
            display_select <= 0;
        end else if (divcnt == HALF_PERIOD - 1) begin
            divcnt <= 0;
            display_select <= ~display_select; // Toggle between displays
        end else begin
            divcnt <= divcnt + 1;            // Increment counter
        end
    end

    // Power multiplexing control for PNP transistors
    assign select0 = display_select;       // Controls PNP for Display 0 (shows s0)
    assign select1 = ~display_select;      // Controls PNP for Display 1 (shows s1), opposite phase

endmodule
